** Profile: "SCHEMATIC1-RC_DC"  [ C:\Cadence\Pspice sim\RC-PSpiceFiles\SCHEMATIC1\RC_DC.sim ] 

** Creating circuit file "RC_DC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\ROG\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 10 1 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\SCHEMATIC1.net" 


.END
