** Profile: "SCHEMATIC1-pp_ac"  [ C:\Cadence\Pspice sim\pp_cascode-PSpiceFiles\SCHEMATIC1\pp_ac.sim ] 

** Creating circuit file "pp_ac.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../pp_cascode-pspicefiles/pp_cascode.lib" 
* From [PSPICE NETLIST] section of C:\Users\ROG\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1Meg 600Meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
