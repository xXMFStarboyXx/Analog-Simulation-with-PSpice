** Profile: "SCHEMATIC1-DC"  [ C:\Cadence\Pspice sim\mycascode-PSpiceFiles\SCHEMATIC1\DC.sim ] 

** Creating circuit file "DC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../mycascode-pspicefiles/mycascode.lib" 
* From [PSPICE NETLIST] section of C:\Users\ROG\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/24.1.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC V_V3 LIST 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
