** Profile: "SCHEMATIC1-tran"  [ C:\Cadence\Pspice sim\smoke_cascode-PSpiceFiles\SCHEMATIC1\tran.sim ] 

** Creating circuit file "tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../smoke_cascode-pspicefiles/smoke_cascode.lib" 
* From [PSPICE NETLIST] section of C:\Users\ROG\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/24.1.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2m 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
