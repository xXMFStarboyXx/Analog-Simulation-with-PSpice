*Wheatstone Bridge
VIN 1 0 10.0VOLT
R1 1 2 2.0ohm
V1 21 2 0
R2 1 3 1ohm
V3 2 22 0
R3 2 0 1ohm
R4 3 0 2ohm
R5 2 3 2ohm
V5 23 2 0
.dc vin 1 2 0.1
.print dc V(VIN) I(r1) I(r2) 
.END