*Wheatstone Bridge
VIN 1 0 10.0VOLT
R1 1 2 2.0ohm
V1 21 2 0
R2 1 3 1ohm
V3 2 22 0
R3 2 0 1ohm
C1 5 3  2pf
R4 4 5 2ohm
C2 0 4  2pf
R5 2 3 2ohm
V5 23 2 0
.END