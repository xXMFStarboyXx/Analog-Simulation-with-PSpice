** Profile: "SCHEMATIC1-bias"  [ C:\Cadence\Pspice sim\digimon-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\Cadence\Pspice sim\digimon-pspicefiles\schematic1\bias\bias_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\ROG\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5 0 
.OPTIONS ADVCONV
.OPTIONS DIGINITSTATE= 0
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
